<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-126.769,11.922,206.052,-206.64</PageViewport>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>29,-14.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>29,-35.5</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>29,-25</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-19.5,3</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>-13.5,3</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-8,3</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>-2.5,3</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_INVERTER</type>
<position>-16.5,-3.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_INVERTER</type>
<position>-10.5,-3.5</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_INVERTER</type>
<position>-5.5,-3.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_INVERTER</type>
<position>0.5,-3.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_OR4</type>
<position>13,-14.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>-19.5,7</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>-13.5,7</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>-8,7</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>-2.5,7</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AE_OR4</type>
<position>13,-25</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>37</ID>
<type>AE_OR4</type>
<position>12.5,-35.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>38</ID>
<type>AE_OR4</type>
<position>12.5,-45.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>40</ID>
<type>AE_OR4</type>
<position>12.5,-56.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>42</ID>
<type>AE_OR4</type>
<position>12.5,-67</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>43</ID>
<type>AE_OR4</type>
<position>12.5,-77.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>12.5,-7.5</position>
<gparam>LABEL_TEXT A0'+A1'+A2'+A3'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>13,-20</position>
<gparam>LABEL_TEXT A0+A1'+A2'+A3'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>12.5,-30</position>
<gparam>LABEL_TEXT A0'+A1+A2'+A3'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>12,-40.5</position>
<gparam>LABEL_TEXT A0+A1+A2'+A3'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>12.5,-50.5</position>
<gparam>LABEL_TEXT A0'+A1'+A2+A3'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>12.5,-61.5</position>
<gparam>LABEL_TEXT A0+A1'+A2+A3'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>12,-72</position>
<gparam>LABEL_TEXT A0'+A1+A2+A3'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AE_OR4</type>
<position>12.5,-88.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>12,-83</position>
<gparam>LABEL_TEXT A0+A1+A2+A3'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AE_OR4</type>
<position>12,-99.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>11.5,-94</position>
<gparam>LABEL_TEXT A0'+A1'+A2'+A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AE_OR4</type>
<position>12,-111</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>11.5,-105.5</position>
<gparam>LABEL_TEXT A0+A1'+A2'+A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>28.5,-45.5</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>28.5,-67</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>28.5,-56.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>28.5,-77.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>28,-88.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>28,-111</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>28,-99.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>34,-14</position>
<gparam>LABEL_TEXT y15</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>33.5,-24.5</position>
<gparam>LABEL_TEXT y14</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>34,-35</position>
<gparam>LABEL_TEXT y13</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>33,-45</position>
<gparam>LABEL_TEXT y12</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>33,-55.5</position>
<gparam>LABEL_TEXT y11</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>33,-66.5</position>
<gparam>LABEL_TEXT y10</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>32.5,-77</position>
<gparam>LABEL_TEXT y9</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>33,-87.5</position>
<gparam>LABEL_TEXT y8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>33.5,-98.5</position>
<gparam>LABEL_TEXT y7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>32.5,-110.5</position>
<gparam>LABEL_TEXT y6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AE_OR4</type>
<position>12.5,-123</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>12,-117.5</position>
<gparam>LABEL_TEXT A0'+A1+A2'+A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>28.5,-123</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>34,-122.5</position>
<gparam>LABEL_TEXT y5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AE_OR4</type>
<position>12.5,-135</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>12,-129.5</position>
<gparam>LABEL_TEXT A0+A1+A2'+A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>28.5,-135</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>33.5,-134.5</position>
<gparam>LABEL_TEXT y4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AE_OR4</type>
<position>12.5,-147</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>12,-141.5</position>
<gparam>LABEL_TEXT A0'+A1'+A2+A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>28.5,-147</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>33.5,-146</position>
<gparam>LABEL_TEXT y3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AE_OR4</type>
<position>13,-159</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>12.5,-153.5</position>
<gparam>LABEL_TEXT A0+A1'+A2+A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>GA_LED</type>
<position>29,-159</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>34,-158</position>
<gparam>LABEL_TEXT y2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AE_OR4</type>
<position>12.5,-170.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>12,-165</position>
<gparam>LABEL_TEXT A0'+A1+A2+A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>GA_LED</type>
<position>28.5,-170.5</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>33.5,-169.5</position>
<gparam>LABEL_TEXT y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AE_OR4</type>
<position>12,-182</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>11.5,-176.5</position>
<gparam>LABEL_TEXT A0+A1+A2+A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>GA_LED</type>
<position>28,-182</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>33,-181</position>
<gparam>LABEL_TEXT y0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>62,-88</position>
<gparam>LABEL_TEXT 4:16 Decoder</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,-179,-19,1</points>
<intersection>-179 35</intersection>
<intersection>-156 38</intersection>
<intersection>-132 29</intersection>
<intersection>-108 23</intersection>
<intersection>-85.5 21</intersection>
<intersection>-64 19</intersection>
<intersection>-42.5 12</intersection>
<intersection>-22 10</intersection>
<intersection>-0.5 3</intersection>
<intersection>1 34</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-19,-0.5,-16.5,-0.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-19,-22,10,-22</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-19,-42.5,9.5,-42.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-19,-64,9.5,-64</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-19,-85.5,9.5,-85.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-19,-108,9,-108</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-19,-132,9.5,-132</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>-19.5,1,-19,1</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>-19,-179,9,-179</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>-19,-156,10,-156</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-181,-13,1</points>
<intersection>-181 37</intersection>
<intersection>-169.5 35</intersection>
<intersection>-134 29</intersection>
<intersection>-122 27</intersection>
<intersection>-87.5 22</intersection>
<intersection>-76.5 20</intersection>
<intersection>-44.5 16</intersection>
<intersection>-34.5 14</intersection>
<intersection>-0.5 7</intersection>
<intersection>1 34</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-13,-0.5,-10.5,-0.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-13,-34.5,9.5,-34.5</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-13,-44.5,9.5,-44.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-13,-76.5,9.5,-76.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-13,-87.5,9.5,-87.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-13,-122,9.5,-122</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-13,-134,9.5,-134</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>-13.5,1,-13,1</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>-13,-169.5,9.5,-169.5</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-13,-181,9,-181</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-183,-7.5,1</points>
<intersection>-183 33</intersection>
<intersection>-171.5 31</intersection>
<intersection>-160 36</intersection>
<intersection>-148 25</intersection>
<intersection>-89.5 20</intersection>
<intersection>-78.5 18</intersection>
<intersection>-68 16</intersection>
<intersection>-57.5 13</intersection>
<intersection>-0.5 4</intersection>
<intersection>1 30</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-7.5,-0.5,-5.5,-0.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-7.5,-57.5,9.5,-57.5</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-7.5,-68,9.5,-68</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-7.5,-78.5,9.5,-78.5</points>
<connection>
<GID>43</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-7.5,-89.5,9.5,-89.5</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-7.5,-148,9.5,-148</points>
<connection>
<GID>84</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-8,1,-7.5,1</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>-7.5,-171.5,9.5,-171.5</points>
<connection>
<GID>104</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>-7.5,-183,9,-183</points>
<connection>
<GID>108</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>-7.5,-160,10,-160</points>
<connection>
<GID>100</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-185,-2,1</points>
<intersection>-185 32</intersection>
<intersection>-173.5 31</intersection>
<intersection>-162 35</intersection>
<intersection>-150 25</intersection>
<intersection>-138 24</intersection>
<intersection>-126 23</intersection>
<intersection>-114 18</intersection>
<intersection>-102.5 16</intersection>
<intersection>-0.5 6</intersection>
<intersection>1 30</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-2,-0.5,0.5,-0.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-2,-102.5,9,-102.5</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-2,-114,9,-114</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-2,-126,9.5,-126</points>
<connection>
<GID>76</GID>
<name>IN_3</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-2,-138,9.5,-138</points>
<connection>
<GID>80</GID>
<name>IN_3</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-2,-150,9.5,-150</points>
<connection>
<GID>84</GID>
<name>IN_3</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-2.5,1,-2,1</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>-2,-173.5,9.5,-173.5</points>
<connection>
<GID>104</GID>
<name>IN_3</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>-2,-185,9,-185</points>
<connection>
<GID>108</GID>
<name>IN_3</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>-2,-162,10,-162</points>
<connection>
<GID>100</GID>
<name>IN_3</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-167.5,-16,-6.5</points>
<intersection>-167.5 35</intersection>
<intersection>-144 28</intersection>
<intersection>-120 26</intersection>
<intersection>-96.5 20</intersection>
<intersection>-74.5 18</intersection>
<intersection>-53.5 16</intersection>
<intersection>-32.5 11</intersection>
<intersection>-11.5 6</intersection>
<intersection>-6.5 33</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-16,-11.5,10,-11.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-16,-32.5,9.5,-32.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-16,-53.5,9.5,-53.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-16,-74.5,9.5,-74.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-16,-96.5,9,-96.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-16,-120,9.5,-120</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-16,-144,9.5,-144</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>-16.5,-6.5,-16,-6.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>-16,-167.5,9.5,-167.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-158,-10,-6.5</points>
<intersection>-158 33</intersection>
<intersection>-146 25</intersection>
<intersection>-110 20</intersection>
<intersection>-98.5 18</intersection>
<intersection>-66 17</intersection>
<intersection>-55.5 14</intersection>
<intersection>-24 11</intersection>
<intersection>-13.5 6</intersection>
<intersection>-6.5 30</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-10,-13.5,10,-13.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-10,-24,10,-24</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-10,-55.5,9.5,-55.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-10,-66,9.5,-66</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-10,-98.5,9,-98.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-10,-110,9,-110</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-10,-146,9.5,-146</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-10.5,-6.5,-10,-6.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>-10,-158,10,-158</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-136,-5,-6.5</points>
<intersection>-136 31</intersection>
<intersection>-124 29</intersection>
<intersection>-112 23</intersection>
<intersection>-100.5 21</intersection>
<intersection>-46.5 16</intersection>
<intersection>-36.5 14</intersection>
<intersection>-26 12</intersection>
<intersection>-15.5 7</intersection>
<intersection>-6.5 36</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-5,-15.5,10,-15.5</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-5,-26,10,-26</points>
<connection>
<GID>36</GID>
<name>IN_2</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-5,-36.5,9.5,-36.5</points>
<connection>
<GID>37</GID>
<name>IN_2</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-5,-46.5,9.5,-46.5</points>
<connection>
<GID>38</GID>
<name>IN_2</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-5,-100.5,9,-100.5</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-5,-112,9,-112</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-5,-124,9.5,-124</points>
<connection>
<GID>76</GID>
<name>IN_2</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>-5,-136,9.5,-136</points>
<connection>
<GID>80</GID>
<name>IN_2</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>-5.5,-6.5,-5,-6.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-91.5,1,-6.5</points>
<intersection>-91.5 17</intersection>
<intersection>-80.5 16</intersection>
<intersection>-70 15</intersection>
<intersection>-59.5 13</intersection>
<intersection>-48.5 10</intersection>
<intersection>-38.5 9</intersection>
<intersection>-28 8</intersection>
<intersection>-17.5 4</intersection>
<intersection>-6.5 26</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1,-17.5,10,-17.5</points>
<connection>
<GID>29</GID>
<name>IN_3</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>1,-28,10,-28</points>
<connection>
<GID>36</GID>
<name>IN_3</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>1,-38.5,9.5,-38.5</points>
<connection>
<GID>37</GID>
<name>IN_3</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>1,-48.5,9.5,-48.5</points>
<connection>
<GID>38</GID>
<name>IN_3</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>1,-59.5,9.5,-59.5</points>
<connection>
<GID>40</GID>
<name>IN_3</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>1,-70,9.5,-70</points>
<connection>
<GID>42</GID>
<name>IN_3</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>1,-80.5,9.5,-80.5</points>
<connection>
<GID>43</GID>
<name>IN_3</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>1,-91.5,9.5,-91.5</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>0.5,-6.5,1,-6.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-14.5,28,-14.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-25,28,-25</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<connection>
<GID>6</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-35.5,28,-35.5</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<connection>
<GID>4</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-45.5,27.5,-45.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>58</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-56.5,27.5,-56.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<connection>
<GID>60</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-67,27.5,-67</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-77.5,27.5,-77.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<connection>
<GID>61</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-88.5,27,-88.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>62</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-99.5,27,-99.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<connection>
<GID>64</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-111,27,-111</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<connection>
<GID>63</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-123,27.5,-123</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>78</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-135,27.5,-135</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<connection>
<GID>82</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-147,27.5,-147</points>
<connection>
<GID>86</GID>
<name>N_in0</name></connection>
<connection>
<GID>84</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-159,28,-159</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<connection>
<GID>102</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-170.5,27.5,-170.5</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-182,27,-182</points>
<connection>
<GID>110</GID>
<name>N_in0</name></connection>
<connection>
<GID>108</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>66.3277,-4.07576,206.737,-96.2822</PageViewport></page 1>
<page 2>
<PageViewport>-68.0104,37.7538,264.81,-180.808</PageViewport></page 2>
<page 3>
<PageViewport>-68.0104,37.7538,264.81,-180.808</PageViewport></page 3>
<page 4>
<PageViewport>-68.0104,37.7538,264.81,-180.808</PageViewport></page 4>
<page 5>
<PageViewport>-68.0104,37.7538,264.81,-180.808</PageViewport></page 5>
<page 6>
<PageViewport>-68.0104,37.7538,264.81,-180.808</PageViewport></page 6>
<page 7>
<PageViewport>-68.0104,37.7538,264.81,-180.808</PageViewport></page 7>
<page 8>
<PageViewport>-68.0104,37.7538,264.81,-180.808</PageViewport></page 8>
<page 9>
<PageViewport>-68.0104,37.7538,264.81,-180.808</PageViewport></page 9></circuit>