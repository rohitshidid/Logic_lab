<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-27.4886,20.3933,90.1302,-56.8464</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-3</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>39.5,-16</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>GA_LED</type>
<position>39.5,-21.5</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-6.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-10.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>-6.5,-2.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>-6.5,-6</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-6.5,-10</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-14.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-6.5,-14</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>44,-15.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>44.5,-10</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>12.5,-36.5</position>
<gparam>LABEL_TEXT Octal To Binary Encoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-18.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-22</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-26</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>-6.5,-18</position>
<gparam>LABEL_TEXT Y4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-6.5,-21.5</position>
<gparam>LABEL_TEXT Y5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>-6.5,-25.5</position>
<gparam>LABEL_TEXT Y6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-30</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>-6.5,-29.5</position>
<gparam>LABEL_TEXT Y7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>39.5,-10.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>44.5,-21</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR4</type>
<position>20.5,-5.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_OR4</type>
<position>20.5,-16</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_OR4</type>
<position>20,-27</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-6.5,8.5,-2.5</points>
<intersection>-6.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-2.5,17.5,-2.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-6.5,8.5,-6.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-15,6.5,-4.5</points>
<intersection>-15 4</intersection>
<intersection>-14.5 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-14.5,6.5,-14.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-4.5,17.5,-4.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>6.5,-15,17.5,-15</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-26,9,-6.5</points>
<intersection>-26 3</intersection>
<intersection>-22 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-22,9,-22</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9,-6.5,17.5,-6.5</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>9,-26,17,-26</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-30,11,-8.5</points>
<intersection>-30 1</intersection>
<intersection>-19 3</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-30,17,-30</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-8.5,17.5,-8.5</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>11,-19,17.5,-19</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-13,8.5,-10.5</points>
<intersection>-13 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-10.5,8.5,-10.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-13,17.5,-13</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-28,4.5,-17</points>
<intersection>-28 4</intersection>
<intersection>-26 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-26,4.5,-26</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-17,17.5,-17</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>4.5,-28,17,-28</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-24,8,-18.5</points>
<intersection>-24 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-18.5,8,-18.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-24,17,-24</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-10.5,33.5,-5.5</points>
<intersection>-10.5 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-10.5,38.5,-10.5</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-5.5,33.5,-5.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-16,38.5,-16</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-27,33.5,-21.5</points>
<intersection>-27 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-21.5,38.5,-21.5</points>
<connection>
<GID>3</GID>
<name>N_in0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-27,33.5,-27</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>12,10.6717,151.4,-80.8717</PageViewport></page 1>
<page 2>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 2>
<page 3>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 3>
<page 4>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 4>
<page 5>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 5>
<page 6>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 6>
<page 7>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 7>
<page 8>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 8>
<page 9>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 9></circuit>