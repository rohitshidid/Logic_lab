<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-27.4886,20.3933,90.1302,-56.8464</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-8,1</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>45,-17</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>GA_LED</type>
<position>45,-22.5</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-8,-2.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>-8,-6.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>-12,1.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>-12,-2</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-12,-6</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>-8,-10.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-12,-10</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>49.5,-16.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>50,-11</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>20,-43.5</position>
<gparam>LABEL_TEXT Decimal To BCD Encoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>-8,-14.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>-8,-18</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>-8,-22</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>-12,-14</position>
<gparam>LABEL_TEXT Y4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-12,-17.5</position>
<gparam>LABEL_TEXT Y5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>-12,-21.5</position>
<gparam>LABEL_TEXT Y6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>-8,-26</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>-12,-25.5</position>
<gparam>LABEL_TEXT Y7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>45,-11.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>50,-22</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>-8,-30</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>-12,-29.5</position>
<gparam>LABEL_TEXT Y8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>-8,-34</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>-12,-33.5</position>
<gparam>LABEL_TEXT Y9</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AE_OR4</type>
<position>16,-5.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_OR4</type>
<position>16,-17</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_OR4</type>
<position>16,-28</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_OR2</type>
<position>28.5,-6.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>45,-27.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>50,-27</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AE_OR2</type>
<position>16,-36</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-2.5,13,-2.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-16,4.5,-4.5</points>
<intersection>-16 3</intersection>
<intersection>-10.5 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-10.5,4.5,-10.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-4.5,13,-4.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>4.5,-16,13,-16</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-27,6,-6.5</points>
<intersection>-27 3</intersection>
<intersection>-18 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-6.5,13,-6.5</points>
<connection>
<GID>28</GID>
<name>IN_2</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6,-18,6,-18</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>6,-27,13,-27</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-31,-0.5,-8.5</points>
<intersection>-31 6</intersection>
<intersection>-26 1</intersection>
<intersection>-20 4</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-26,-0.5,-26</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-8.5,13,-8.5</points>
<connection>
<GID>28</GID>
<name>IN_3</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-0.5,-20,13,-20</points>
<connection>
<GID>29</GID>
<name>IN_3</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-0.5,-31,13,-31</points>
<connection>
<GID>30</GID>
<name>IN_3</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-14,3.5,-6.5</points>
<intersection>-14 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-6.5,3.5,-6.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-14,13,-14</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-29,7,-18</points>
<intersection>-29 3</intersection>
<intersection>-22 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-22,7,-22</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-18,13,-18</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>7,-29,13,-29</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-25,3.5,-14.5</points>
<intersection>-25 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-14.5,3.5,-14.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-25,13,-25</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-5.5,25.5,-5.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-11.5,37.5,-6.5</points>
<intersection>-11.5 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-11.5,44,-11.5</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-6.5,37.5,-6.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-37,-2.5,-12</points>
<intersection>-37 6</intersection>
<intersection>-34 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-34,-2.5,-34</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2.5,-12,19.5,-12</points>
<intersection>-2.5 0</intersection>
<intersection>19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19.5,-12,19.5,-7.5</points>
<intersection>-12 2</intersection>
<intersection>-7.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19.5,-7.5,25.5,-7.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>19.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-2.5,-37,13,-37</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>-2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-17,44,-17</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-28,32,-22.5</points>
<intersection>-28 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-22.5,44,-22.5</points>
<connection>
<GID>3</GID>
<name>N_in0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-28,32,-28</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-35,3.5,-30</points>
<intersection>-35 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-30,3.5,-30</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-35,13,-35</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-36,34,-27.5</points>
<intersection>-36 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-27.5,44,-27.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-36,34,-36</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>12,10.6717,151.4,-80.8717</PageViewport></page 1>
<page 2>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 2>
<page 3>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 3>
<page 4>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 4>
<page 5>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 5>
<page 6>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 6>
<page 7>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 7>
<page 8>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 8>
<page 9>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 9></circuit>