<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-52.0537,45.635,188.104,-112.075</PageViewport>
<gate>
<ID>2</ID>
<type>AM_MUX_16x1</type>
<position>72,-19.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_10</ID>6 </input>
<input>
<ID>IN_11</ID>5 </input>
<input>
<ID>IN_12</ID>4 </input>
<input>
<ID>IN_13</ID>3 </input>
<input>
<ID>IN_14</ID>2 </input>
<input>
<ID>IN_15</ID>1 </input>
<input>
<ID>IN_2</ID>14 </input>
<input>
<ID>IN_3</ID>13 </input>
<input>
<ID>IN_4</ID>12 </input>
<input>
<ID>IN_5</ID>11 </input>
<input>
<ID>IN_6</ID>10 </input>
<input>
<ID>IN_7</ID>9 </input>
<input>
<ID>IN_8</ID>8 </input>
<input>
<ID>IN_9</ID>7 </input>
<output>
<ID>OUT</ID>33 </output>
<input>
<ID>SEL_0</ID>39 </input>
<input>
<ID>SEL_1</ID>38 </input>
<input>
<ID>SEL_2</ID>37 </input>
<input>
<ID>SEL_3</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>4</ID>
<type>AM_MUX_16x1</type>
<position>72,-50</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<input>
<ID>IN_10</ID>22 </input>
<input>
<ID>IN_11</ID>21 </input>
<input>
<ID>IN_12</ID>20 </input>
<input>
<ID>IN_13</ID>19 </input>
<input>
<ID>IN_14</ID>18 </input>
<input>
<ID>IN_15</ID>17 </input>
<input>
<ID>IN_2</ID>30 </input>
<input>
<ID>IN_3</ID>29 </input>
<input>
<ID>IN_4</ID>28 </input>
<input>
<ID>IN_5</ID>27 </input>
<input>
<ID>IN_6</ID>26 </input>
<input>
<ID>IN_7</ID>25 </input>
<input>
<ID>IN_8</ID>24 </input>
<input>
<ID>IN_9</ID>23 </input>
<output>
<ID>OUT</ID>34 </output>
<input>
<ID>SEL_0</ID>39 </input>
<input>
<ID>SEL_1</ID>38 </input>
<input>
<ID>SEL_2</ID>37 </input>
<input>
<ID>SEL_3</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>27,-1.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>27,-3.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>27,-5.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>27,-7.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>27,-9.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>27,-11.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>27,-13.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>27,-15.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>27,-17.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>27,-19.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>27,-21.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>27,-23.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>27,-25.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>27,-27.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>27,-29.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>27,-31.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>27,-35</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>27,-37</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>27,-39</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>27,-41</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>27,-43</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>27,-45</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>27,-47</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>27,-49</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>27,-51</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>27,-53</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>27,-55</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>27,-57</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>27,-59</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>27,-61</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>27,-63</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>27,-65</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_OR2</type>
<position>105.5,-31</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>GA_LED</type>
<position>112.5,-31</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>69,-2.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>75,-2.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>79,-2.5</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>72,-2.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>24,-1.5</position>
<gparam>LABEL_TEXT D31</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>24,-3.5</position>
<gparam>LABEL_TEXT D30</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>24,-5.5</position>
<gparam>LABEL_TEXT D29</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>24,-7.5</position>
<gparam>LABEL_TEXT D28</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>24,-9.5</position>
<gparam>LABEL_TEXT D27</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>24,-11.5</position>
<gparam>LABEL_TEXT D26</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>24,-13.5</position>
<gparam>LABEL_TEXT D25</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>24,-15.5</position>
<gparam>LABEL_TEXT D24</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>24,-17</position>
<gparam>LABEL_TEXT D23</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>24,-19</position>
<gparam>LABEL_TEXT D22</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>24,-21</position>
<gparam>LABEL_TEXT D21</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>24,-23</position>
<gparam>LABEL_TEXT D20</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>24,-25</position>
<gparam>LABEL_TEXT D19</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>24,-27</position>
<gparam>LABEL_TEXT D18</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>24,-29</position>
<gparam>LABEL_TEXT D17</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>24,-31</position>
<gparam>LABEL_TEXT D16</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>24,-34.5</position>
<gparam>LABEL_TEXT D15</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>24,-36.5</position>
<gparam>LABEL_TEXT D14</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>24,-38.5</position>
<gparam>LABEL_TEXT D13</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>24,-40.5</position>
<gparam>LABEL_TEXT D12</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>24,-42.5</position>
<gparam>LABEL_TEXT D11</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>24,-44.5</position>
<gparam>LABEL_TEXT D10</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>24,-46.5</position>
<gparam>LABEL_TEXT D9</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>24,-48.5</position>
<gparam>LABEL_TEXT D8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>24,-50.5</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>24,-52.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>24,-54.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>24,-56.5</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>24,-58.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>24,-60.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>24.5,-62.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>24,-64.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>69,-0.5</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>72,-0.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>75,-0.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>79,-0.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-12,58.5,-1.5</points>
<intersection>-12 1</intersection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-12,69,-12</points>
<connection>
<GID>2</GID>
<name>IN_15</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-1.5,58.5,-1.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-13,57.5,-3.5</points>
<intersection>-13 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-13,69,-13</points>
<connection>
<GID>2</GID>
<name>IN_14</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-3.5,57.5,-3.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-14,56.5,-5.5</points>
<intersection>-14 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-14,69,-14</points>
<connection>
<GID>2</GID>
<name>IN_13</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-5.5,56.5,-5.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-15,55.5,-7.5</points>
<intersection>-15 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-15,69,-15</points>
<connection>
<GID>2</GID>
<name>IN_12</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-7.5,55.5,-7.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-16,54.5,-9.5</points>
<intersection>-16 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-16,69,-16</points>
<connection>
<GID>2</GID>
<name>IN_11</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-9.5,54.5,-9.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-17,53.5,-11.5</points>
<intersection>-17 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-17,69,-17</points>
<connection>
<GID>2</GID>
<name>IN_10</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-11.5,53.5,-11.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-18,53,-13.5</points>
<intersection>-18 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-18,69,-18</points>
<connection>
<GID>2</GID>
<name>IN_9</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-13.5,53,-13.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-19,52,-15.5</points>
<intersection>-19 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-19,69,-19</points>
<connection>
<GID>2</GID>
<name>IN_8</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-15.5,52,-15.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-20,51,-17.5</points>
<intersection>-20 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-20,69,-20</points>
<connection>
<GID>2</GID>
<name>IN_7</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-17.5,51,-17.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-21,50,-19.5</points>
<intersection>-21 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-21,69,-21</points>
<connection>
<GID>2</GID>
<name>IN_6</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-19.5,50,-19.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-22,49,-21.5</points>
<intersection>-22 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-22,69,-22</points>
<connection>
<GID>2</GID>
<name>IN_5</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-21.5,49,-21.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-23.5,49,-23</points>
<intersection>-23.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-23,69,-23</points>
<connection>
<GID>2</GID>
<name>IN_4</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-23.5,49,-23.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-25.5,49,-24</points>
<intersection>-25.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-24,69,-24</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-25.5,49,-25.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-27.5,49.5,-25</points>
<intersection>-27.5 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-25,69,-25</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-27.5,49.5,-27.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-29.5,50.5,-26</points>
<intersection>-29.5 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-26,69,-26</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-29.5,50.5,-29.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-31.5,51.5,-27</points>
<intersection>-31.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-27,69,-27</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-31.5,51.5,-31.5</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-42.5,61.5,-35</points>
<intersection>-42.5 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-42.5,69,-42.5</points>
<connection>
<GID>4</GID>
<name>IN_15</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-35,61.5,-35</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-43.5,60.5,-37</points>
<intersection>-43.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-43.5,69,-43.5</points>
<connection>
<GID>4</GID>
<name>IN_14</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-37,60.5,-37</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-44.5,59.5,-39</points>
<intersection>-44.5 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-44.5,69,-44.5</points>
<connection>
<GID>4</GID>
<name>IN_13</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-39,59.5,-39</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-45.5,58.5,-41</points>
<intersection>-45.5 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-45.5,69,-45.5</points>
<connection>
<GID>4</GID>
<name>IN_12</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-41,58.5,-41</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-46.5,57.5,-43</points>
<intersection>-46.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-46.5,69,-46.5</points>
<connection>
<GID>4</GID>
<name>IN_11</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-43,57.5,-43</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-47.5,56.5,-45</points>
<intersection>-47.5 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-47.5,69,-47.5</points>
<connection>
<GID>4</GID>
<name>IN_10</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-45,56.5,-45</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-48.5,55.5,-47</points>
<intersection>-48.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-48.5,69,-48.5</points>
<connection>
<GID>4</GID>
<name>IN_9</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-47,55.5,-47</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-49.5,54.5,-49</points>
<intersection>-49.5 1</intersection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-49.5,69,-49.5</points>
<connection>
<GID>4</GID>
<name>IN_8</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-49,54.5,-49</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-51,49,-50.5</points>
<intersection>-51 2</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-50.5,69,-50.5</points>
<connection>
<GID>4</GID>
<name>IN_7</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-51,49,-51</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-53,49,-51.5</points>
<intersection>-53 2</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-51.5,69,-51.5</points>
<connection>
<GID>4</GID>
<name>IN_6</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-53,49,-53</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-55,49.5,-52.5</points>
<intersection>-55 2</intersection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-52.5,69,-52.5</points>
<connection>
<GID>4</GID>
<name>IN_5</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-55,49.5,-55</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-57,50.5,-53.5</points>
<intersection>-57 2</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-53.5,69,-53.5</points>
<connection>
<GID>4</GID>
<name>IN_4</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-57,50.5,-57</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-59,51.5,-54.5</points>
<intersection>-59 2</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-54.5,69,-54.5</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-59,51.5,-59</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-61,52.5,-55.5</points>
<intersection>-61 2</intersection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-55.5,69,-55.5</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-61,52.5,-61</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-63,53.5,-56.5</points>
<intersection>-63 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-56.5,69,-56.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-63,53.5,-63</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-65,54.5,-57.5</points>
<intersection>-65 2</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-57.5,69,-57.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-65,54.5,-65</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-30,88.5,-19.5</points>
<intersection>-30 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-30,102.5,-30</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-19.5,88.5,-19.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-50,88.5,-32</points>
<intersection>-50 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-32,102.5,-32</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-50,88.5,-50</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108.5,-31,111.5,-31</points>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<connection>
<GID>39</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-37,76,-7.5</points>
<intersection>-37 4</intersection>
<intersection>-10 5</intersection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>69,-7.5,69,-4.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-7.5,76,-7.5</points>
<intersection>69 1</intersection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>70.5,-37,76,-37</points>
<intersection>70.5 6</intersection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>70.5,-10,76,-10</points>
<connection>
<GID>2</GID>
<name>SEL_3</name></connection>
<intersection>76 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>70.5,-40.5,70.5,-37</points>
<connection>
<GID>4</GID>
<name>SEL_3</name></connection>
<intersection>-37 4</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-38.5,77,-7</points>
<intersection>-38.5 4</intersection>
<intersection>-10 5</intersection>
<intersection>-7 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>72,-7,72,-4.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>72,-7,77,-7</points>
<intersection>72 1</intersection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>71.5,-38.5,77,-38.5</points>
<intersection>71.5 6</intersection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>71.5,-10,77,-10</points>
<connection>
<GID>2</GID>
<name>SEL_2</name></connection>
<intersection>77 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>71.5,-40.5,71.5,-38.5</points>
<connection>
<GID>4</GID>
<name>SEL_2</name></connection>
<intersection>-38.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-39.5,78.5,-6.5</points>
<intersection>-39.5 4</intersection>
<intersection>-10 5</intersection>
<intersection>-6.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>75,-6.5,75,-4.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75,-6.5,78.5,-6.5</points>
<intersection>75 1</intersection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>72.5,-39.5,78.5,-39.5</points>
<intersection>72.5 6</intersection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>72.5,-10,78.5,-10</points>
<connection>
<GID>2</GID>
<name>SEL_1</name></connection>
<intersection>78.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>72.5,-40.5,72.5,-39.5</points>
<connection>
<GID>4</GID>
<name>SEL_1</name></connection>
<intersection>-39.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-40.5,79.5,-6</points>
<intersection>-40.5 5</intersection>
<intersection>-10 6</intersection>
<intersection>-6 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>79,-6,79,-4.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>79,-6,79.5,-6</points>
<intersection>79 1</intersection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>73.5,-40.5,79.5,-40.5</points>
<connection>
<GID>4</GID>
<name>SEL_0</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>73.5,-10,79.5,-10</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>146.78,-24.7703,292.866,-120.704</PageViewport></page 1>
<page 2>
<PageViewport>0,71.4106,439.646,-217.303</PageViewport></page 2>
<page 3>
<PageViewport>0,71.4106,439.646,-217.303</PageViewport></page 3>
<page 4>
<PageViewport>164.867,-36.6221,274.779,-108.8</PageViewport></page 4>
<page 5>
<PageViewport>0,71.4106,439.646,-217.303</PageViewport></page 5>
<page 6>
<PageViewport>0,71.4106,439.646,-217.303</PageViewport></page 6>
<page 7>
<PageViewport>0,71.4106,439.646,-217.303</PageViewport></page 7>
<page 8>
<PageViewport>0,71.4106,439.646,-217.303</PageViewport></page 8>
<page 9>
<PageViewport>0,71.4106,439.646,-217.303</PageViewport></page 9></circuit>