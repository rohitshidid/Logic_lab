<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-214.92,143.211,277.561,-180.198</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-73,17.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>-42.5,6</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>GA_LED</type>
<position>-42.5,0.5</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-73,14</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>-73,10</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>-77,18</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>-77,14.5</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-77,10.5</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>-73,6</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-77,6.5</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>-38,6.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>-37.5,12</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>-62.5,-16</position>
<gparam>LABEL_TEXT 8:3 Encoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>-73,2</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>-73,-1.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>-73,-5.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>-77,2.5</position>
<gparam>LABEL_TEXT Y4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-77,-1</position>
<gparam>LABEL_TEXT Y5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>-77,-5</position>
<gparam>LABEL_TEXT Y6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>-73,-9.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>-77,-9</position>
<gparam>LABEL_TEXT Y7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>-42.5,11.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>-37.5,1</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR4</type>
<position>-56.5,14.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_OR4</type>
<position>-56.5,5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_OR4</type>
<position>-56.5,-5.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,14,-65.5,17.5</points>
<intersection>14 2</intersection>
<intersection>17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65.5,17.5,-59.5,17.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71,14,-65.5,14</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,6,-64.5,15.5</points>
<intersection>6 2</intersection>
<intersection>15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,15.5,-59.5,15.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71,6,-59.5,6</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-4.5,-66.5,13.5</points>
<intersection>-4.5 3</intersection>
<intersection>-1.5 2</intersection>
<intersection>13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66.5,13.5,-59.5,13.5</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71,-1.5,-66.5,-1.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-66.5,-4.5,-59.5,-4.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,-9.5,-63.5,11.5</points>
<intersection>-9.5 2</intersection>
<intersection>-8.5 4</intersection>
<intersection>2 3</intersection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,11.5,-59.5,11.5</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71,-9.5,-63.5,-9.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-63.5,2,-59.5,2</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-63.5,-8.5,-59.5,-8.5</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>-63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68.5,8,-59.5,8</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-68.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-68.5,8,-68.5,10</points>
<intersection>8 1</intersection>
<intersection>10 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-71,10,-68.5,10</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-68.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-6.5,-64.5,4</points>
<intersection>-6.5 3</intersection>
<intersection>-5.5 1</intersection>
<intersection>4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71,-5.5,-64.5,-5.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-64.5,4,-59.5,4</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-64.5,-6.5,-59.5,-6.5</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,-2.5,-68.5,2</points>
<intersection>-2.5 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71,2,-68.5,2</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-68.5,-2.5,-59.5,-2.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,11.5,-48,14.5</points>
<intersection>11.5 1</intersection>
<intersection>14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48,11.5,-43.5,11.5</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>-48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,14.5,-48,14.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>-48 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,5,-48,6</points>
<intersection>5 2</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48,6,-43.5,6</points>
<connection>
<GID>2</GID>
<name>N_in0</name></connection>
<intersection>-48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,5,-48,5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>-48 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,-5.5,-48,0.5</points>
<intersection>-5.5 2</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48,0.5,-43.5,0.5</points>
<connection>
<GID>3</GID>
<name>N_in0</name></connection>
<intersection>-48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-5.5,-48,-5.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-48 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>12,10.6717,151.4,-80.8717</PageViewport></page 1>
<page 2>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 2>
<page 3>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 3>
<page 4>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 4>
<page 5>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 5>
<page 6>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 6>
<page 7>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 7>
<page 8>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 8>
<page 9>
<PageViewport>0,10.6717,139.4,-80.8717</PageViewport></page 9></circuit>